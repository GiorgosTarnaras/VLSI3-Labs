library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity led_mux is
    port (
        clk     : in  std_logic;
        reset   : in  std_logic;  
        in0     : in  std_logic_vector(7 downto 0);
        in1     : in  std_logic_vector(7 downto 0);
        in2     : in  std_logic_vector(7 downto 0);
        in3     : in  std_logic_vector(7 downto 0);
        an      : out std_logic_vector(3 downto 0);  
        sseg    : out std_logic_vector(7 downto 0)
    );
end led_mux;

architecture arch of led_mux is

    signal counter : unsigned(15 downto 0);
    signal display_sel : unsigned(1 downto 0);
    
begin
	process(clk, reset)
    begin
        if reset = '1' then
            counter <= (others => '0');
        elsif rising_edge(clk) then
            counter <= counter + 1;
        end if;
    end process;

    display_sel <= std_logic_vector(counter(15 downto 14));
    
    with display_sel select
        sseg <= in0 when "00",
                in1 when "01",
                in2 when "10",
                in3 when others;
    
    with display_sel select
        an <= "1110" when "00",  
              "1101" when "01",  
              "1011" when "10",  
              "0111" when others; 

end arch;
